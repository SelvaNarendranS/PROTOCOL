VCD info: dumpfile dump.vcd opened for output.

Time = 0 | rst = 0 | data_in = 0(00000000) | tx = 1 | busy = 0 |rx = x | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 0 | rxst = 0
Time = 1000 | rst = 0 | data_in = 0(00000000) | tx = 1 | busy = 0 |rx = 1 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 0 | rxst = 0
Time = 100000 | rst = 1 | data_in = 0(00000000) | tx = 1 | busy = 0 |rx = 1 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 0 | rxst = 0

------------------------- Sending Data:  40 | parity en & type  = 1 & EVEN-----------------------
Time = 105000 | rst = 1 | data_in = 40(00101000) | tx = 1 | busy = 1 |rx = 1 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 1 | rxst = 0
Time = 104265000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 1 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 0
Time = 104266000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 0
Time = 110610000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 1
Time = 162610000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 520905000 | rst = 1 | data_in = 40(00101000) | tx = 1 | busy = 1 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 520906000 | rst = 1 | data_in = 40(00101000) | tx = 1 | busy = 1 |rx = 1 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 625065000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 1 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 625066000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 729225000 | rst = 1 | data_in = 40(00101000) | tx = 1 | busy = 1 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 729226000 | rst = 1 | data_in = 40(00101000) | tx = 1 | busy = 1 |rx = 1 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 833385000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 1 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 833386000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 937545000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 3 | rxst = 2
Time = 994610000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 3 | rxst = 3
Time = 1041705000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 4 | rxst = 3
Time = 1098610000 | rst = 1 | data_in = 40(00101000) | tx = 0 | busy = 1 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 4 | rxst = 4
Time = 1145865000 | rst = 1 | data_in = 40(00101000) | tx = 1 | busy = 0 |rx = 0 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 0 | rxst = 4
Time = 1145866000 | rst = 1 | data_in = 40(00101000) | tx = 1 | busy = 0 |rx = 1 | data_out = 0(00000000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 0 | rxst = 4
Time = 1202610000 | rst = 1 | data_in = 40(00101000) | tx = 1 | busy = 0 |rx = 1 | data_out = 40(00101000) | done = 1 | frm_err = 0 | pty_err = 0 | txst = 0 | rxst = 0
	------------------------------------------------------------
			 SUCCESS: Received  40 correctly
	--------------------------------------------------------------

------------------------- Sending Data:  85 | parity en & type  = 1 & ODD-----------------------
Time = 1202915000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 1 | frm_err = 0 | pty_err = 0 | txst = 1 | rxst = 0
Time = 1209110000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 1 | rxst = 0
Time = 1250025000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 0
Time = 1250026000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 0
Time = 1254610000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 1
Time = 1306610000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1354185000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1354186000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1458345000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1458346000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1562505000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1562506000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1666665000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1666666000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1770825000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1770826000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1874985000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1874986000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1979145000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 1979146000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 2083305000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 3 | rxst = 2
Time = 2083306000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 3 | rxst = 2
Time = 2138610000 | rst = 1 | data_in = 85(01010101) | tx = 0 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 3 | rxst = 3
Time = 2187465000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 0 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 4 | rxst = 3
Time = 2187466000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 4 | rxst = 3
Time = 2242610000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 1 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 4 | rxst = 4
Time = 2291625000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 0 |rx = 1 | data_out = 40(00101000) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 0 | rxst = 4
Time = 2346610000 | rst = 1 | data_in = 85(01010101) | tx = 1 | busy = 0 |rx = 1 | data_out = 85(01010101) | done = 1 | frm_err = 0 | pty_err = 0 | txst = 0 | rxst = 0
	------------------------------------------------------------
			 SUCCESS: Received  85 correctly
	--------------------------------------------------------------

------------------------- Sending Data: 123 | parity en & type  = 0 & ODD-----------------------
Time = 2346915000 | rst = 1 | data_in = 123(01111011) | tx = 1 | busy = 1 |rx = 1 | data_out = 85(01010101) | done = 1 | frm_err = 0 | pty_err = 0 | txst = 1 | rxst = 0
Time = 2353110000 | rst = 1 | data_in = 123(01111011) | tx = 1 | busy = 1 |rx = 1 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 1 | rxst = 0
Time = 2395785000 | rst = 1 | data_in = 123(01111011) | tx = 0 | busy = 1 |rx = 1 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 0
Time = 2395786000 | rst = 1 | data_in = 123(01111011) | tx = 0 | busy = 1 |rx = 0 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 0
Time = 2398610000 | rst = 1 | data_in = 123(01111011) | tx = 0 | busy = 1 |rx = 0 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 1
Time = 2450610000 | rst = 1 | data_in = 123(01111011) | tx = 0 | busy = 1 |rx = 0 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 2499945000 | rst = 1 | data_in = 123(01111011) | tx = 1 | busy = 1 |rx = 0 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 2499946000 | rst = 1 | data_in = 123(01111011) | tx = 1 | busy = 1 |rx = 1 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 2708265000 | rst = 1 | data_in = 123(01111011) | tx = 0 | busy = 1 |rx = 1 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 2708266000 | rst = 1 | data_in = 123(01111011) | tx = 0 | busy = 1 |rx = 0 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 2812425000 | rst = 1 | data_in = 123(01111011) | tx = 1 | busy = 1 |rx = 0 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 2812426000 | rst = 1 | data_in = 123(01111011) | tx = 1 | busy = 1 |rx = 1 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 2 | rxst = 2
Time = 3229065000 | rst = 1 | data_in = 123(01111011) | tx = 0 | busy = 1 |rx = 1 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 4 | rxst = 2
Time = 3229066000 | rst = 1 | data_in = 123(01111011) | tx = 0 | busy = 1 |rx = 0 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 4 | rxst = 2
Time = 3282610000 | rst = 1 | data_in = 123(01111011) | tx = 0 | busy = 1 |rx = 0 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 4 | rxst = 4
Time = 3333225000 | rst = 1 | data_in = 123(01111011) | tx = 1 | busy = 0 |rx = 0 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 0 | rxst = 4
Time = 3333226000 | rst = 1 | data_in = 123(01111011) | tx = 1 | busy = 0 |rx = 1 | data_out = 85(01010101) | done = 0 | frm_err = 0 | pty_err = 0 | txst = 0 | rxst = 4
Time = 3386610000 | rst = 1 | data_in = 123(01111011) | tx = 1 | busy = 0 |rx = 1 | data_out = 123(01111011) | done = 1 | frm_err = 0 | pty_err = 0 | txst = 0 | rxst = 0
	------------------------------------------------------------
			 SUCCESS: Received 123 correctly
	--------------------------------------------------------------

testbench.v:94: $finish called at 3387910000 (1ps)